magic
tech scmos
timestamp 1702426510
<< nwell >>
rect -132 30 -113 31
rect -132 -5 190 30
<< ntransistor >>
rect -103 -65 -100 -56
rect -61 -65 -58 -56
rect -45 -65 -42 -56
rect -29 -65 -26 -56
rect 3 -65 6 -56
rect 19 -65 22 -56
rect 37 -65 40 -56
rect 51 -65 54 -56
rect 64 -65 67 -56
rect 82 -65 85 -56
rect 105 -65 108 -56
rect 120 -65 123 -56
rect 131 -65 134 -56
rect 161 -65 164 -56
<< ptransistor >>
rect -103 1 -100 8
rect -61 1 -58 8
rect -45 1 -42 8
rect -29 1 -26 8
rect 3 1 6 8
rect 19 1 22 8
rect 37 1 40 8
rect 51 1 54 8
rect 64 1 67 8
rect 82 1 85 8
rect 105 1 108 8
rect 120 1 123 8
rect 131 1 134 8
rect 161 1 164 8
<< ndiffusion >>
rect -118 -64 -113 -56
rect -108 -64 -103 -56
rect -118 -65 -103 -64
rect -100 -57 -61 -56
rect -100 -65 -98 -57
rect -92 -59 -61 -57
rect -92 -63 -72 -59
rect -68 -63 -61 -59
rect -92 -65 -61 -63
rect -58 -60 -45 -56
rect -58 -65 -55 -60
rect -50 -65 -45 -60
rect -42 -59 -29 -56
rect -42 -63 -37 -59
rect -33 -63 -29 -59
rect -42 -65 -29 -63
rect -26 -65 -15 -56
rect -10 -65 3 -56
rect 6 -65 19 -56
rect 22 -59 37 -56
rect 22 -65 26 -59
rect 32 -65 37 -59
rect 40 -62 43 -56
rect 49 -62 51 -56
rect 40 -65 51 -62
rect 54 -60 64 -56
rect 54 -65 56 -60
rect 62 -65 64 -60
rect 67 -63 71 -56
rect 76 -63 82 -56
rect 67 -65 82 -63
rect 85 -63 91 -56
rect 96 -63 105 -56
rect 85 -65 105 -63
rect 108 -65 120 -56
rect 123 -65 131 -56
rect 134 -58 161 -56
rect 134 -65 144 -58
rect 153 -65 161 -58
rect 164 -62 170 -56
rect 176 -62 187 -56
rect 164 -65 187 -62
<< pdiffusion >>
rect -121 6 -103 8
rect -121 1 -113 6
rect -108 1 -103 6
rect -100 1 -98 8
rect -92 1 -91 8
rect -88 6 -61 8
rect -88 2 -76 6
rect -72 2 -61 6
rect -88 1 -61 2
rect -58 4 -55 8
rect -50 4 -45 8
rect -58 1 -45 4
rect -42 6 -29 8
rect -42 2 -39 6
rect -35 2 -29 6
rect -42 1 -29 2
rect -26 1 -15 8
rect -10 1 3 8
rect 6 1 19 8
rect 22 3 28 8
rect 34 3 37 8
rect 22 1 37 3
rect 40 6 51 8
rect 40 1 43 6
rect 49 1 51 6
rect 54 4 56 8
rect 61 4 64 8
rect 54 1 64 4
rect 67 6 82 8
rect 67 1 72 6
rect 77 1 82 6
rect 85 7 105 8
rect 85 1 91 7
rect 96 1 105 7
rect 108 1 120 8
rect 123 1 131 8
rect 134 3 137 8
rect 144 3 147 8
rect 134 1 147 3
rect 151 1 153 8
rect 158 1 161 8
rect 164 6 181 8
rect 164 1 170 6
rect 176 1 181 6
<< ndcontact >>
rect -113 -64 -108 -56
rect -98 -65 -92 -57
rect -72 -63 -68 -59
rect -55 -65 -50 -60
rect -37 -63 -33 -59
rect -15 -65 -10 -56
rect 26 -65 32 -59
rect 43 -62 49 -56
rect 56 -65 62 -60
rect 71 -63 76 -56
rect 91 -63 96 -56
rect 144 -65 153 -58
rect 170 -62 176 -56
<< pdcontact >>
rect -113 1 -108 6
rect -98 1 -92 8
rect -76 2 -72 6
rect -55 4 -50 8
rect -39 2 -35 6
rect -15 1 -10 8
rect 28 3 34 8
rect 43 1 49 6
rect 56 4 61 8
rect 72 1 77 6
rect 91 1 96 7
rect 137 3 144 8
rect 153 1 158 8
rect 170 1 176 6
<< psubstratepcontact >>
rect -72 -97 156 -88
<< nsubstratencontact >>
rect -75 21 145 25
<< polysilicon >>
rect -103 8 -100 12
rect -61 8 -58 12
rect -45 8 -42 12
rect -29 8 -26 12
rect 3 8 6 12
rect 19 8 22 12
rect 37 8 40 12
rect 51 8 54 12
rect 64 8 67 13
rect 82 8 85 13
rect 105 8 108 13
rect 120 8 123 13
rect 131 8 134 13
rect 161 8 164 12
rect -103 -15 -100 1
rect -61 -7 -58 1
rect -103 -56 -100 -20
rect -61 -56 -58 -11
rect -45 -29 -42 1
rect -45 -56 -42 -33
rect -29 -37 -26 1
rect 3 -7 6 1
rect -29 -56 -26 -41
rect 3 -56 6 -11
rect 19 -33 22 1
rect 37 -7 40 1
rect 19 -56 22 -37
rect 37 -56 40 -11
rect 51 -33 54 1
rect 51 -56 54 -37
rect 64 -42 67 1
rect 82 -25 85 1
rect 105 -7 108 1
rect 64 -56 67 -46
rect 82 -56 85 -29
rect 105 -56 108 -11
rect 120 -27 123 1
rect 120 -56 123 -31
rect 131 -42 134 1
rect 161 -15 164 1
rect 131 -56 134 -46
rect 161 -56 164 -20
rect -103 -70 -100 -65
rect -61 -70 -58 -65
rect -45 -70 -42 -65
rect -29 -70 -26 -65
rect 3 -70 6 -65
rect 19 -70 22 -65
rect 37 -70 40 -65
rect 51 -70 54 -65
rect 64 -70 67 -65
rect 82 -70 85 -65
rect 105 -70 108 -65
rect 120 -70 123 -65
rect 131 -70 134 -65
rect 161 -71 164 -65
<< polycontact >>
rect -63 -11 -58 -7
rect -103 -20 -97 -15
rect -47 -33 -42 -29
rect 1 -11 6 -7
rect -31 -41 -26 -37
rect 35 -11 40 -7
rect 17 -37 22 -33
rect 49 -37 54 -33
rect 103 -11 108 -7
rect 79 -29 85 -25
rect 64 -46 71 -42
rect 119 -31 123 -27
rect 158 -20 164 -15
rect 128 -46 134 -42
<< metal1 >>
rect -108 21 -75 25
rect 145 21 170 25
rect -129 11 -101 15
rect -113 -14 -108 1
rect -105 -7 -101 11
rect -98 8 -92 21
rect -55 8 -50 21
rect -24 11 -3 15
rect -76 1 -72 2
rect -39 1 -35 2
rect -76 -3 -35 1
rect -24 -7 -20 11
rect -105 -11 -63 -7
rect -58 -11 -20 -7
rect -128 -20 -108 -14
rect -15 -15 -10 1
rect -6 -7 -3 11
rect 28 8 34 21
rect 56 8 61 21
rect 82 12 103 16
rect 43 -4 77 1
rect 82 -7 86 12
rect -6 -11 1 -7
rect 6 -11 35 -7
rect 40 -11 86 -7
rect -97 -20 -10 -15
rect -129 -33 -126 -27
rect -113 -56 -108 -20
rect -15 -25 -10 -20
rect 91 -15 96 1
rect 99 -11 103 12
rect 137 8 144 21
rect 153 8 158 21
rect 91 -20 158 -15
rect -15 -29 79 -25
rect -91 -33 -47 -29
rect -42 -33 -18 -29
rect -105 -41 -31 -37
rect -105 -70 -101 -41
rect -72 -56 -33 -52
rect -126 -76 -101 -70
rect -72 -59 -68 -56
rect -37 -59 -33 -56
rect -98 -88 -92 -65
rect -55 -88 -50 -65
rect -30 -78 -26 -41
rect -22 -69 -18 -33
rect -15 -56 -10 -29
rect 8 -37 17 -33
rect 22 -37 49 -33
rect 54 -37 88 -33
rect 8 -69 12 -37
rect -22 -73 12 -69
rect 16 -46 64 -42
rect 71 -46 82 -42
rect 16 -78 20 -46
rect 43 -56 76 -51
rect -30 -82 20 -78
rect 26 -88 32 -65
rect 56 -88 62 -65
rect 79 -78 82 -46
rect 85 -70 88 -37
rect 91 -56 96 -20
rect 170 -22 176 1
rect 115 -70 119 -27
rect 170 -28 180 -22
rect 85 -74 119 -70
rect 126 -46 128 -42
rect 126 -78 130 -46
rect 170 -56 176 -28
rect 79 -82 130 -78
rect 144 -88 153 -65
rect -104 -97 -72 -88
rect 156 -97 189 -88
<< m2contact >>
rect -126 -33 -119 -27
rect -99 -33 -91 -27
<< metal2 >>
rect -119 -33 -99 -27
<< labels >>
rlabel metal1 -78 -94 -78 -94 1 Gnd
rlabel metal1 -85 22 -85 22 1 Vdd
rlabel m2contact -98 -31 -98 -31 3 B
rlabel metal1 -96 -39 -96 -39 3 C
rlabel metal1 178 -25 178 -25 1 Sum
rlabel metal1 -117 -17 -117 -17 1 Cout
rlabel metal1 -96 -10 -96 -10 3 A
<< end >>
