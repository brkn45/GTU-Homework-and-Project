magic
tech scmos
timestamp 1703957753
<< metal1 >>
rect -3 71 1 76
rect 98 63 135 67
rect -25 35 16 39
rect -25 1 -20 35
rect 101 20 106 26
rect 113 21 117 31
rect 131 21 135 63
rect 101 16 109 20
rect -34 -4 -20 1
rect -25 -56 -20 -4
rect -11 9 16 13
rect 104 11 109 16
rect -11 -47 -7 9
rect 104 7 118 11
rect 6 0 12 5
rect 93 0 135 4
rect -4 -24 2 -19
rect 93 -28 98 0
rect 114 -10 124 -6
rect -25 -60 6 -56
rect 106 -67 111 -11
rect 219 -21 223 -17
rect 118 -42 124 -22
rect 118 -43 126 -42
rect 118 -45 127 -43
rect -11 -81 -5 -70
rect 104 -71 111 -67
rect -11 -82 18 -81
rect 161 -82 166 -32
rect -11 -86 14 -82
rect 99 -86 166 -82
rect 6 -95 8 -90
<< m2contact >>
rect 113 16 118 21
rect 118 7 123 12
rect 106 -11 111 -6
rect -11 -53 -4 -47
rect -11 -70 -3 -64
rect 118 -22 124 -16
<< metal2 >>
rect 106 16 113 20
rect 106 -6 111 16
rect 118 -16 123 7
rect -11 -64 -5 -53
use 2mux  2mux_2
timestamp 1703881869
transform 1 0 181 0 1 1
box -68 -46 41 30
use 2mux  2mux_1
timestamp 1703881869
transform 1 0 67 0 1 -49
box -68 -46 41 30
use 2mux  2mux_0
timestamp 1703881869
transform 1 0 68 0 1 46
box -68 -46 41 30
<< labels >>
rlabel metal1 96 -3 96 -3 1 Vdd4
rlabel metal1 219 -21 223 -17 7 Y4
rlabel metal1 -31 -2 -31 -2 3 s0
rlabel metal1 -2 74 -2 74 5 d1b
rlabel metal1 7 2 7 2 1 d0b
rlabel metal1 -3 -22 -3 -21 1 d3b
rlabel metal1 7 -93 7 -93 1 d2b
rlabel metal1 115 -8 115 -8 1 s1
rlabel metal1 122 -84 122 -84 1 Gnd4
<< end >>
