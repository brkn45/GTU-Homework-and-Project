magic
tech scmos
timestamp 1703881869
<< nwell >>
rect -66 -4 41 25
<< ntransistor >>
rect -45 -29 -43 -25
rect -24 -29 -22 -25
rect -11 -29 -9 -25
rect 4 -29 6 -25
rect 18 -29 20 -25
<< ptransistor >>
rect -45 3 -43 7
rect -24 3 -22 7
rect -11 3 -9 7
rect 4 3 6 7
rect 18 3 20 7
<< ndiffusion >>
rect -46 -29 -45 -25
rect -43 -29 -40 -25
rect -36 -29 -33 -25
rect -30 -29 -29 -25
rect -25 -29 -24 -25
rect -22 -29 -11 -25
rect -9 -29 -5 -25
rect -1 -29 4 -25
rect 6 -29 18 -25
rect 20 -29 23 -25
rect 27 -29 32 -25
<< pdiffusion >>
rect -52 3 -50 7
rect -46 3 -45 7
rect -43 3 -40 7
rect -36 3 -35 7
rect -32 3 -30 7
rect -26 3 -24 7
rect -22 3 -19 7
rect -15 3 -11 7
rect -9 3 -4 7
rect 0 3 4 7
rect 6 3 10 7
rect 14 3 18 7
rect 20 3 24 7
rect 28 3 35 7
<< ndcontact >>
rect -50 -29 -46 -25
rect -40 -29 -36 -25
rect -29 -29 -25 -25
rect -5 -29 -1 -25
rect 23 -29 27 -25
<< pdcontact >>
rect -50 3 -46 7
rect -40 3 -36 7
rect -30 3 -26 7
rect -19 3 -15 7
rect -4 3 0 7
rect 10 3 14 7
rect 24 3 28 7
<< psubstratepcontact >>
rect -51 -37 -47 -33
rect -43 -37 -38 -33
rect -34 -37 -25 -33
rect -12 -37 -7 -33
rect 0 -37 5 -33
rect 9 -37 13 -33
rect 18 -37 23 -33
rect 28 -37 32 -33
<< nsubstratencontact >>
rect -50 17 -46 21
rect -38 17 -33 21
rect -22 17 -17 21
rect -1 17 4 21
rect 25 17 29 21
<< polysilicon >>
rect -60 25 20 27
rect -45 14 -9 16
rect -45 7 -43 14
rect -24 7 -22 10
rect -11 7 -9 14
rect 4 7 6 10
rect 18 7 20 25
rect -45 -7 -43 3
rect -44 -11 -43 -7
rect -45 -25 -43 -11
rect -24 -25 -22 3
rect -11 -25 -9 3
rect 4 -7 6 3
rect 5 -11 6 -7
rect 4 -25 6 -11
rect 18 -25 20 3
rect -45 -32 -43 -29
rect -24 -41 -22 -29
rect -11 -32 -9 -29
rect 4 -32 6 -29
rect 18 -32 20 -29
rect -51 -43 -22 -41
<< polycontact >>
rect -64 25 -60 30
rect -48 -11 -44 -7
rect 1 -11 5 -7
rect -55 -46 -51 -41
<< metal1 >>
rect -68 25 -64 30
rect -46 17 -38 21
rect -33 17 -22 21
rect -17 17 -1 21
rect 4 17 25 21
rect 29 17 31 21
rect -50 7 -46 17
rect -19 7 -15 17
rect -40 -7 -36 3
rect -4 10 28 14
rect -4 7 0 10
rect 24 7 28 10
rect -30 0 -26 3
rect -4 0 0 3
rect -30 -4 0 0
rect -61 -11 -48 -7
rect -40 -11 1 -7
rect -40 -25 -36 -11
rect 10 -18 14 3
rect -5 -22 38 -18
rect -5 -25 -1 -22
rect -50 -33 -46 -29
rect -29 -33 -25 -29
rect 23 -33 27 -29
rect -53 -37 -51 -33
rect -47 -37 -43 -33
rect -38 -37 -34 -33
rect -25 -37 -12 -33
rect -7 -37 0 -33
rect 5 -37 9 -33
rect 13 -37 18 -33
rect 23 -37 28 -33
rect -59 -46 -55 -41
<< labels >>
rlabel metal1 -60 -9 -60 -9 1 s
rlabel metal1 -58 -44 -58 -44 1 d0
rlabel metal1 -67 27 -67 27 4 d1
rlabel nsubstratencontact -47 19 -47 19 1 vdd
rlabel nsubstratencontact -47 19 -47 19 1 Vdd
rlabel psubstratepcontact -50 -35 -50 -35 1 Gnd
rlabel metal1 36 -20 36 -20 7 Y
<< end >>
