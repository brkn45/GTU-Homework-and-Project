magic
tech scmos
timestamp 1699462543
<< nwell >>
rect -16 -2 12 27
<< ntransistor >>
rect -3 -17 -1 -13
<< ptransistor >>
rect -3 6 -1 10
<< ndiffusion >>
rect -5 -17 -3 -13
rect -1 -17 1 -13
rect 5 -17 6 -13
<< pdiffusion >>
rect -9 6 -8 10
rect -4 6 -3 10
rect -1 6 1 10
rect 5 6 6 10
<< ndcontact >>
rect -9 -17 -5 -13
rect 1 -17 5 -13
<< pdcontact >>
rect -8 6 -4 10
rect 1 6 5 10
<< nsubstratencontact >>
rect -12 19 -8 23
rect -2 19 2 23
rect -9 -32 -5 -28
rect 0 -32 4 -28
<< polysilicon >>
rect -3 10 -1 13
rect -3 -4 -1 6
rect -2 -8 -1 -4
rect -3 -13 -1 -8
rect -3 -22 -1 -17
<< polycontact >>
rect -7 -8 -2 -4
<< metal1 >>
rect -13 19 -12 23
rect -8 19 -2 23
rect 2 19 6 23
rect -13 18 6 19
rect -8 10 -4 18
rect -11 -8 -7 -4
rect 1 -5 5 6
rect 1 -10 10 -5
rect 1 -13 5 -10
rect -9 -27 -5 -17
rect -9 -28 5 -27
rect -5 -32 0 -28
rect 4 -32 5 -28
<< labels >>
rlabel metal1 -3 -29 -3 -29 1 gnd!
rlabel metal1 -6 21 -6 21 1 vdd!
rlabel metal1 -11 -6 -11 -6 3 in!
rlabel metal1 10 -8 10 -8 7 out
<< end >>
